library verilog;
use verilog.vl_types.all;
entity add4_sv_unit is
end add4_sv_unit;
