library verilog;
use verilog.vl_types.all;
entity mdr_decoder_sv_unit is
end mdr_decoder_sv_unit;
